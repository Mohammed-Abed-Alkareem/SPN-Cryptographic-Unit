package spn_tb_pkg;
    
    import uvm_pkg::*;
    import spn_cu_pkg::*;
    
    `include "spn_seq_item.sv"
    `include "spn_sequencer.sv"
    `include "spn_sequence.sv"
    `include "spn_driver.sv"
    `include "spn_monitor.sv"
    `include "spn_scoreboard.sv"
    `include "spn_agent.sv"
    `include "spn_env.sv"
    `include "spn_base_test.sv"
    `include "spn_test.sv"
    `include "spn_test_encrypt.sv"
    `include "spn_test_decrypt.sv"
endpackage